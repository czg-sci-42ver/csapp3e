// `include "E4.13.1.v"
module moduleName (
    ports
);
    input ports;
    wire clock;
endmodule

// always #1 clock = ~clock;
